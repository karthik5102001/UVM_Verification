package pack;

  import uvm_pkg::*;

`include "uvm_macros.svh"

`include "Transaction.sv"
`include "sequence_1.sv"
`include "Driver.sv"
`include "Monitor_1.sv"
`include "Agent_1.sv"
`include "Scoreboard.sv"
`include "Env.sv"
`include "Test.sv"

endpackage